`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 14.10.2019 21:59:04
// Design Name: 
// Module Name: mux32to1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux32to1(
    output Y,
    input [31:0] A,
    input [4:0] C
    );
    wire [31:0] Y1;
    assign #1 Y1[0]=A[0]&~C[0]&~C[1]&~C[2]&~C[3]&~C[4];
    assign #1 Y1[1]=A[1]&C[0]&~C[1]&~C[2]&~C[3]&~C[4];
    assign #1 Y1[2]=A[2]&~C[0]&C[1]&~C[2]&~C[3]&~C[4];
    assign #1 Y1[3]=A[3]&C[0]&C[1]&~C[2]&~C[3]&~C[4];
    assign #1 Y1[4]=A[4]&~C[0]&~C[1]&C[2]&~C[3]&~C[4];
    assign #1 Y1[5]=A[5]&C[0]&~C[1]&C[2]&~C[3]&~C[4];
    assign #1 Y1[6]=A[6]&~C[0]&C[1]&C[2]&~C[3]&~C[4];
    assign #1 Y1[7]=A[7]&C[0]&C[1]&C[2]&~C[3]&~C[4];
    assign #1 Y1[8]=A[8]&~C[0]&~C[1]&~C[2]&C[3]&~C[4];
    assign #1 Y1[9]=A[9]&C[0]&~C[1]&~C[2]&C[3]&~C[4];
    assign #1 Y1[10]=A[10]&~C[0]&C[1]&~C[2]&C[3]&~C[4];
    assign #1 Y1[11]=A[11]&C[0]&C[1]&~C[2]&C[3]&~C[4];
    assign #1 Y1[12]=A[12]&~C[0]&~C[1]&C[2]&C[3]&~C[4];
    assign #1 Y1[13]=A[13]&C[0]&~C[1]&C[2]&C[3]&~C[4];
    assign #1 Y1[14]=A[14]&~C[0]&C[1]&C[2]&C[3]&~C[4];
    assign #1 Y1[15]=A[15]&C[0]&C[1]&C[2]&C[3]&~C[4];
    assign #1 Y1[16]=A[16]&~C[0]&~C[1]&~C[2]&~C[3]&C[4];
    assign #1 Y1[17]=A[17]&C[0]&~C[1]&~C[2]&~C[3]&C[4];
    assign #1 Y1[18]=A[18]&~C[0]&C[1]&~C[2]&~C[3]&C[4];
    assign #1 Y1[19]=A[19]&C[0]&C[1]&~C[2]&~C[3]&C[4];
    assign #1 Y1[20]=A[20]&~C[0]&~C[1]&C[2]&~C[3]&C[4];
    assign #1 Y1[21]=A[21]&C[0]&~C[1]&C[2]&~C[3]&C[4];
    assign #1 Y1[22]=A[22]&~C[0]&C[1]&C[2]&~C[3]&C[4];
    assign #1 Y1[23]=A[23]&C[0]&C[1]&C[2]&~C[3]&C[4];
    assign #1 Y1[24]=A[24]&~C[0]&~C[1]&~C[2]&C[3]&C[4];
    assign #1 Y1[25]=A[25]&C[0]&~C[1]&~C[2]&C[3]&C[4];
    assign #1 Y1[26]=A[26]&~C[0]&C[1]&~C[2]&C[3]&C[4];
    assign #1 Y1[27]=A[27]&C[0]&C[1]&~C[2]&C[3]&C[4];
    assign #1 Y1[28]=A[28]&~C[0]&~C[1]&C[2]&C[3]&C[4];
    assign #1 Y1[29]=A[29]&C[0]&~C[1]&C[2]&C[3]&C[4];
    assign #1 Y1[30]=A[30]&~C[0]&C[1]&C[2]&C[3]&C[4];
    assign #1 Y1[31]=A[31]&C[0]&C[1]&C[2]&C[3]&C[4];
    assign #1 Y=Y1[0]|Y1[1]|Y1[2]|Y1[3]|Y1[4]|Y1[5]|Y1[6]|Y1[7]|Y1[8]|Y1[9]|Y1[10]|Y1[11]|Y1[12]|Y1[13]|Y1[14]|Y1[15]|Y1[16]|Y1[17]|Y1[18]|Y1[19]|Y1[20]|Y1[21]|Y1[22]|Y1[23]|Y1[24]|Y1[25]|Y1[26]|Y1[27]|Y1[28]|Y1[29]|Y1[30]|Y1[31];
endmodule
