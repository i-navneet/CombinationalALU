`timescale 1ns/1ps
//delay for OR/AND gate-1ns NOT delay is 0
//////////////////////////////////////////////////////////////////////////////////
// Company: Indian Institute of Technology
// Engineer: Navtejpreet Singh
//            Navneet Kumar
// 
// Create Date: 16.10.2019 00:28:32
// Design Name: 
// Module Name: CLA4bit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module CLA4bit(
    output [3:0] S,
    output C,
    output C1,
    input[3:0] A,
    input[3:0] B,
    input Cin
);
//wire P and G saves carry propagate and carry generation
// carry wires save carry for inwards sum
//P[i]=A[i]|B[i] G[i]=A[i]&B[i]
//Sum is generated by these carry
wire [3:0] P,G;
wire [3:0]Carry;
    assign #1 P[0]=A[0]|B[0];
    assign #1 G[0]=A[0]&B[0];
    assign #2 S[0] = A[0] ^ B[0] ^ Cin;
    assign #2 Carry[1] = A[0] & B[0] | A[0] & Cin | B[0] & Cin;

    assign #1 P[1]=A[1]|B[1];
    assign #1 G[1]=A[1]&B[1];
    assign #2 S[1] = A[1] ^ B[1] ^ Carry[1];
    assign #2 Carry[2] = A[1] & B[1] | A[1] & Carry[1] | B[1] & Carry[1];

    assign #1 P[2]=A[2]|B[2];
    assign #1 G[2]=A[2]&B[2];
    assign #2 S[2] = A[2] ^ B[2] ^ Carry[2];
    assign #2 Carry[3] = A[2] & B[2] | A[2] & Carry[2] | B[2] & Carry[2];

    assign #1 P[3]=A[3]|B[3];
    assign #1 G[3]=A[3]&B[3];
    assign #2 S[3]=A[3] ^ B[3] ^ Carry[3];
//Carry is given by G|P&Cin
assign #2 C = G[0]&P[1]&P[2]&P[3] | G[1]&P[2]&P[3] | G[2]&P[3]| G[3] | P[0]&P[1]&P[2]&P[3]&Cin;
//C1 is second last carry
assign #2 C1 = G[2] | G[1]&P[2] | G[0]&P[1]&P[2] | P[0]&P[1]&P[2]&Cin; 
endmodule